library ieee;
use ieee.std_logic_1164.all;

package types is
	subtype tGameBoard is std_logic_vector(0 to 159);
	

end package types;