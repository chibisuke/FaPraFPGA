library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package constants is
	constant COEFF_LEN_MAX: integer := 1000;

	type tCoeff is array(0 to COEFF_LEN_MAX-1) of signed(23 downto 0);
	type tCoeffArr is array(0 to 3) of tCoeff;
	subtype tCoeffLenRange is integer range 0 to 1000;
	type tCoeffLen is array(0 to 3) of tCoeffLenRange;
	
	constant COEFFICIENTS_1_LEN: integer range 0 to COEFF_LEN_MAX := 129;
	constant COEFFICIENTS_1: tCoeff := (
		x"000078",x"0000a5",x"0000d7",x"00010d",x"000146",x"000180",x"0001b8",x"0001ed",
		x"00021a",x"00023e",x"000256",x"00025e",x"000253",x"000234",x"0001fd",x"0001ad",
		x"000142",x"0000bc",x"00001b",x"ffff5f",x"fffe89",x"fffd9d",x"fffc9d",x"fffb8f",
		x"fffa76",x"fff95b",x"fff843",x"fff736",x"fff63d",x"fff560",x"fff4aa",x"fff422",
		x"fff3d2",x"fff3c4",x"fff400",x"fff48e",x"fff574",x"fff6b9",x"fff861",x"fffa70",
		x"fffce7",x"ffffc5",x"000309",x"0006b1",x"000ab5",x"000f0e",x"0013b4",x"00189a",
		x"001db5",x"0022f6",x"00284e",x"002dae",x"003304",x"00383f",x"003d4e",x"004220",
		x"0046a3",x"004ac9",x"004e82",x"0051c1",x"00547a",x"0056a2",x"005833",x"005926",
		x"005977",x"005926",x"005833",x"0056a2",x"00547a",x"0051c1",x"004e82",x"004ac9",
		x"0046a3",x"004220",x"003d4e",x"00383f",x"003304",x"002dae",x"00284e",x"0022f6",
		x"001db5",x"00189a",x"0013b4",x"000f0e",x"000ab5",x"0006b1",x"000309",x"ffffc5",
		x"fffce7",x"fffa70",x"fff861",x"fff6b9",x"fff574",x"fff48e",x"fff400",x"fff3c4",
		x"fff3d2",x"fff422",x"fff4aa",x"fff560",x"fff63d",x"fff736",x"fff843",x"fff95b",
		x"fffa76",x"fffb8f",x"fffc9d",x"fffd9d",x"fffe89",x"ffff5f",x"00001b",x"0000bc",
		x"000142",x"0001ad",x"0001fd",x"000234",x"000253",x"00025e",x"000256",x"00023e",
		x"00021a",x"0001ed",x"0001b8",x"000180",x"000146",x"00010d",x"0000d7",x"0000a5",
		x"000078",
		others=>x"000000"	
	);
	
	constant COEFFICIENTS_2_LEN: integer range 0 to 1000 := 129;
	constant COEFFICIENTS_2: tCoeff := (
		x"ffff90",x"ffff60",x"ffff30",x"ffff00",x"fffec0",x"fffe80",x"fffe50",x"fffe20",
		x"fffdf0",x"fffdd0",x"fffdb0",x"fffdb0",x"fffdb0",x"fffdd0",x"fffe10",x"fffe60",
		x"fffec0",x"ffff50",x"fffff0",x"0000a0",x"000170",x"000260",x"000360",x"000470",
		x"000580",x"0006a0",x"0007b0",x"0008c0",x"0009c0",x"000a90",x"000b50",x"000bd0",
		x"000c20",x"000c30",x"000bf0",x"000b60",x"000a80",x"000940",x"000790",x"000580",
		x"000310",x"000030",x"fffd00",x"fff960",x"fff550",x"fff100",x"ffec60",x"ffe770",
		x"ffe260",x"ffdd20",x"ffd7c0",x"ffd270",x"ffcd10",x"ffc7e0",x"ffc2d0",x"ffbe00",
		x"ffb980",x"ffb550",x"ffb1a0",x"ffae60",x"ffabb0",x"ffa980",x"ffa7f0",x"ffa700",
		x"07a700",x"ffa700",x"ffa7f0",x"ffa980",x"ffabb0",x"ffae60",x"ffb1a0",x"ffb550",
		x"ffb980",x"ffbe00",x"ffc2d0",x"ffc7e0",x"ffcd10",x"ffd270",x"ffd7c0",x"ffdd20",
		x"ffe260",x"ffe770",x"ffec60",x"fff100",x"fff550",x"fff960",x"fffd00",x"000030",
		x"000310",x"000580",x"000790",x"000940",x"000a80",x"000b60",x"000bf0",x"000c30",
		x"000c20",x"000bd0",x"000b50",x"000a90",x"0009c0",x"0008c0",x"0007b0",x"0006a0",
		x"000580",x"000470",x"000360",x"000260",x"000170",x"0000a0",x"fffff0",x"ffff50",
		x"fffec0",x"fffe60",x"fffe10",x"fffdd0",x"fffdb0",x"fffdb0",x"fffdb0",x"fffdd0",
		x"fffdf0",x"fffe20",x"fffe50",x"fffe80",x"fffec0",x"ffff00",x"ffff30",x"ffff60",
		x"ffff90",
		others=>x"000000"
	);
	
	constant COEFFICIENTS_3_LEN: integer range 0 to 1000 := 129;
	constant COEFFICIENTS_3: tCoeff := (
		x"001E2F",x"FFF66D",x"FFF6EB",x"FFF6DD",x"FFF66E",x"FFF5C4",x"FFF4FE",x"FFF43B",
		x"FFF396",x"FFF325",x"FFF2FD",x"FFF32E",x"FFF3C6",x"FFF4CB",x"FFF644",x"FFF82F",
		x"FFFA84",x"FFFD39",x"00003F",x"000382",x"0006E8",x"000A54",x"000DAD",x"0010D2",
		x"0013A1",x"001602",x"0017D4",x"001901",x"001975",x"001921",x"0017FE",x"001609",
		x"00134A",x"000FCD",x"000BA0",x"0006F8",x"0001C5",x"FFFC5C",x"FFF6DB",x"FFF162",
		x"FFEC23",x"FFE74F",x"FFE315",x"FFDF9B",x"FFDD01",x"FFDB63",x"FFDAD3",x"FFDB5F",
		x"FFDD0B",x"FFDFCF",x"FFE39B",x"FFE855",x"FFEDDB",x"FFF407",x"FFFAA9",x"00018B",
		x"000876",x"000F36",x"001597",x"001B5B",x"00205E",x"00246F",x"002770",x"002948",
		x"0029E7",x"002948",x"002770",x"00246F",x"00205E",x"001B5B",x"001597",x"000F36",
		x"000876",x"00018B",x"FFFAA9",x"FFF407",x"FFEDDB",x"FFE855",x"FFE39B",x"FFDFCF",
		x"FFDD0B",x"FFDB5F",x"FFDAD3",x"FFDB63",x"FFDD01",x"FFDF9B",x"FFE315",x"FFE74F",
		x"FFEC23",x"FFF162",x"FFF6DB",x"FFFC5C",x"0001C5",x"0006F8",x"000BA0",x"000FCD",
		x"00134A",x"001609",x"0017FE",x"001921",x"001975",x"001901",x"0017D4",x"001602",
		x"0013A1",x"0010D2",x"000DAD",x"000A54",x"0006E8",x"000382",x"00003F",x"FFFD39",
		x"FFFA84",x"FFF82F",x"FFF644",x"FFF4CB",x"FFF3C6",x"FFF32E",x"FFF2FD",x"FFF325",
		x"FFF396",x"FFF43B",x"FFF4FE",x"FFF5C4",x"FFF66E",x"FFF6DD",x"FFF6EB",x"FFF66D",
		x"001E2F",
		others=>x"000000"
	);
	
	constant COEFFICIENTS_4_LEN: integer range 0 to 1000 := 129;
	constant COEFFICIENTS_4: tCoeff := (
		x"FFF8BA",x"FFF944",x"FFFA16",x"FFFB20",x"FFFC50",x"FFFD90",x"FFFEC9",x"FFFFE3",
		x"0000C8",x"000164",x"0001A3",x"000177",x"0000D7",x"FFFFBD",x"FFFE2C",x"FFFC29",
		x"FFF9C2",x"FFF70A",x"FFF41A",x"FFF10F",x"FFEE09",x"FFEB2C",x"FFE89D",x"FFE680",
		x"FFE4F9",x"FFE426",x"FFE424",x"FFE508",x"FFE6E0",x"FFE9B3",x"FFED7F",x"FFF239",
		x"FFF7CD",x"FFFE1E",x"000506",x"000C59",x"0013E4",x"001B70",x"0022C2",x"00299E",
		x"002FCA",x"00350E",x"003936",x"003C16",x"003D8A",x"003D76",x"003BCC",x"003887",
		x"0033B1",x"002D5E",x"0025AE",x"001CCE",x"0012F4",x"00085E",x"FFFD52",x"FFF21A",
		x"FFE704",x"FFDC5C",x"FFD26E",x"FFC980",x"FFC1D3",x"FFBB9D",x"FFB70C",x"FFB441",
		x"083894",x"FFB441",x"FFB70C",x"FFBB9D",x"FFC1D3",x"FFC980",x"FFD26E",x"FFDC5C",
		x"FFE704",x"FFF21A",x"FFFD52",x"00085E",x"0012F4",x"001CCE",x"0025AE",x"002D5E",
		x"0033B1",x"003887",x"003BCC",x"003D76",x"003D8A",x"003C16",x"003936",x"00350E",
		x"002FCA",x"00299E",x"0022C2",x"001B70",x"0013E4",x"000C59",x"000506",x"FFFE1E",
		x"FFF7CD",x"FFF239",x"FFED7F",x"FFE9B3",x"FFE6E0",x"FFE508",x"FFE424",x"FFE426",
		x"FFE4F9",x"FFE680",x"FFE89D",x"FFEB2C",x"FFEE09",x"FFF10F",x"FFF41A",x"FFF70A",
		x"FFF9C2",x"FFFC29",x"FFFE2C",x"FFFFBD",x"0000D7",x"000177",x"0001A3",x"000164",
		x"0000C8",x"FFFFE3",x"FFFEC9",x"FFFD90",x"FFFC50",x"FFFB20",x"FFFA16",x"FFF944",
		x"FFF8BA",
		others=>x"000000"
	);
	
	
	constant COEFFICIENTS_5_LEN: integer range 0 to 1000 := 999;
	constant COEFFICIENTS_5: tCoeff := (
		x"fffe56",x"0001bb",x"000136",x"0000f4",x"0000d7",x"0000ce",x"0000d0",x"0000d8" ,
		x"0000e2",x"0000ed",x"0000f9",x"000103",x"00010d",x"000115",x"00011b",x"000120" ,
		x"000122",x"000123",x"000121",x"00011d",x"000117",x"00010e",x"000104",x"0000f7" ,
		x"0000e9",x"0000d8",x"0000c7",x"0000b3",x"00009f",x"000089",x"000073",x"00005c" ,
		x"000046",x"00002f",x"000018",x"000003",x"ffffee",x"ffffda",x"ffffc8",x"ffffb7" ,
		x"ffffa8",x"ffff9b",x"ffff91",x"ffff88",x"ffff82",x"ffff7f",x"ffff7d",x"ffff7e" ,
		x"ffff82",x"ffff87",x"ffff8f",x"ffff99",x"ffffa4",x"ffffb1",x"ffffbf",x"ffffce" ,
		x"ffffde",x"ffffee",x"ffffff",x"00000f",x"00001f",x"00002e",x"00003d",x"00004a" ,
		x"000056",x"000060",x"000068",x"00006e",x"000072",x"000074",x"000074",x"000072" ,
		x"00006d",x"000067",x"00005f",x"000054",x"000049",x"00003c",x"00002d",x"00001e" ,
		x"00000e",x"fffffe",x"ffffee",x"ffffdf",x"ffffcf",x"ffffc1",x"ffffb4",x"ffffa8" ,
		x"ffff9e",x"ffff95",x"ffff8e",x"ffff8a",x"ffff87",x"ffff87",x"ffff8a",x"ffff8d" ,
		x"ffff95",x"ffff9c",x"ffffa7",x"ffffb4",x"ffffc1",x"ffffd0",x"ffffe0",x"fffff1" ,
		x"000001",x"000012",x"000024",x"000034",x"000044",x"000052",x"00005f",x"00006a" ,
		x"000074",x"00007c",x"000081",x"000084",x"000084",x"000082",x"00007e",x"000077" ,
		x"00006f",x"000063",x"000056",x"000048",x"000037",x"000026",x"000014",x"000001" ,
		x"ffffee",x"ffffdb",x"ffffc9",x"ffffb7",x"ffffa7",x"ffff98",x"ffff8b",x"ffff80" ,
		x"ffff77",x"ffff71",x"ffff6d",x"ffff6c",x"ffff6e",x"ffff72",x"ffff79",x"ffff82" ,
		x"ffff8e",x"ffff9d",x"ffffad",x"ffffbe",x"ffffd2",x"ffffe6",x"fffffb",x"000010" ,
		x"000025",x"00003a",x"00004e",x"000060",x"000071",x"000080",x"00008d",x"000098" ,
		x"0000a0",x"0000a5",x"0000a7",x"0000a5",x"0000a1",x"00009a",x"000090",x"000083" ,
		x"000074",x"000062",x"00004f",x"00003a",x"000023",x"00000c",x"fffff4",x"ffffdc" ,
		x"ffffc4",x"ffffae",x"ffff98",x"ffff84",x"ffff73",x"ffff63",x"ffff57",x"ffff4d" ,
		x"ffff47",x"ffff44",x"ffff44",x"ffff48",x"ffff4f",x"ffff5a",x"ffff67",x"ffff78" ,
		x"ffff8b",x"ffffa1",x"ffffb9",x"ffffd2",x"ffffec",x"000007",x"000022",x"00003d" ,
		x"000057",x"000070",x"000087",x"00009b",x"0000ad",x"0000bc",x"0000c8",x"0000d0" ,
		x"0000d5",x"0000d6",x"0000d2",x"0000cb",x"0000c0",x"0000b2",x"0000a0",x"00008a" ,
		x"000073",x"000058",x"00003c",x"00001e",x"000000",x"ffffe1",x"ffffc2",x"ffffa5" ,
		x"ffff88",x"ffff6e",x"ffff55",x"ffff40",x"ffff2e",x"ffff1f",x"ffff15",x"ffff0f" ,
		x"ffff0d",x"ffff0f",x"ffff16",x"ffff21",x"ffff31",x"ffff44",x"ffff5c",x"ffff76" ,
		x"ffff93",x"ffffb3",x"ffffd4",x"fffff7",x"00001a",x"00003d",x"00005f",x"000080" ,
		x"0000a0",x"0000bc",x"0000d5",x"0000eb",x"0000fd",x"00010a",x"000112",x"000116" ,
		x"000114",x"00010e",x"000102",x"0000f2",x"0000dd",x"0000c3",x"0000a6",x"000085" ,
		x"000062",x"00003c",x"000015",x"ffffed",x"ffffc4",x"ffff9d",x"ffff76",x"ffff52" ,
		x"ffff31",x"ffff13",x"fffef8",x"fffee3",x"fffed2",x"fffec7",x"fffec1",x"fffec1" ,
		x"fffec7",x"fffed3",x"fffee5",x"fffefb",x"ffff17",x"ffff38",x"ffff5d",x"ffff85" ,
		x"ffffaf",x"ffffdc",x"00000a",x"000039",x"000067",x"000093",x"0000be",x"0000e6" ,
		x"000109",x"000129",x"000143",x"000158",x"000167",x"00016f",x"000171",x"00016c" ,
		x"000160",x"00014e",x"000135",x"000116",x"0000f2",x"0000c9",x"00009b",x"00006b" ,
		x"000037",x"000002",x"ffffcc",x"ffff96",x"ffff62",x"ffff2f",x"ffff00",x"fffed5" ,
		x"fffeaf",x"fffe8e",x"fffe74",x"fffe61",x"fffe55",x"fffe51",x"fffe54",x"fffe60" ,
		x"fffe73",x"fffe8e",x"fffeb0",x"fffed9",x"ffff08",x"ffff3c",x"ffff74",x"ffffb0" ,
		x"ffffee",x"00002d",x"00006d",x"0000ab",x"0000e7",x"000120",x"000155",x"000184" ,
		x"0001ac",x"0001cd",x"0001e6",x"0001f7",x"0001ff",x"0001fd",x"0001f2",x"0001de" ,
		x"0001c1",x"00019a",x"00016c",x"000136",x"0000fa",x"0000b8",x"000072",x"000028" ,
		x"ffffdd",x"ffff91",x"ffff45",x"fffefc",x"fffeb7",x"fffe76",x"fffe3b",x"fffe08" ,
		x"fffddd",x"fffdbc",x"fffda5",x"fffd98",x"fffd96",x"fffda0",x"fffdb5",x"fffdd6" ,
		x"fffe01",x"fffe36",x"fffe75",x"fffebc",x"ffff0b",x"ffff5f",x"ffffb8",x"000014" ,
		x"000072",x"0000cf",x"00012a",x"000181",x"0001d3",x"00021e",x"000260",x"000299" ,
		x"0002c7",x"0002e8",x"0002fc",x"000303",x"0002fb",x"0002e5",x"0002c1",x"000290" ,
		x"000251",x"000206",x"0001af",x"00014f",x"0000e6",x"000077",x"000003",x"ffff8d" ,
		x"ffff15",x"fffe9f",x"fffe2d",x"fffdc1",x"fffd5d",x"fffd03",x"fffcb4",x"fffc74" ,
		x"fffc42",x"fffc21",x"fffc12",x"fffc14",x"fffc2a",x"fffc52",x"fffc8c",x"fffcd9" ,
		x"fffd36",x"fffda4",x"fffe20",x"fffea8",x"ffff3a",x"ffffd5",x"000075",x"000118" ,
		x"0001ba",x"000259",x"0002f3",x"000383",x"000407",x"00047d",x"0004e1",x"000531" ,
		x"00056c",x"00058e",x"000598",x"000587",x"00055b",x"000515",x"0004b3",x"000437" ,
		x"0003a2",x"0002f5",x"000234",x"00015f",x"00007b",x"ffff8a",x"fffe91",x"fffd93" ,
		x"fffc95",x"fffb9b",x"fffaaa",x"fff9c6",x"fff8f4",x"fff838",x"fff798",x"fff717" ,
		x"fff6ba",x"fff684",x"fff678",x"fff699",x"fff6ea",x"fff76d",x"fff821",x"fff909" ,
		x"fffa24",x"fffb71",x"fffcef",x"fffe9d",x"000076",x"000278",x"00049f",x"0006e7" ,
		x"00094b",x"000bc5",x"000e4f",x"0010e4",x"00137c",x"001612",x"00189f",x"001b1d" ,
		x"001d83",x"001fce",x"0021f5",x"0023f3",x"0025c4",x"002761",x"0028c6",x"0029f0" ,
		x"002adc",x"002b85",x"002bec",x"002c0f",x"002bec",x"002b85",x"002adc",x"0029f0" ,
		x"0028c6",x"002761",x"0025c4",x"0023f3",x"0021f5",x"001fce",x"001d83",x"001b1d" ,
		x"00189f",x"001612",x"00137c",x"0010e4",x"000e4f",x"000bc5",x"00094b",x"0006e7" ,
		x"00049f",x"000278",x"000076",x"fffe9d",x"fffcef",x"fffb71",x"fffa24",x"fff909" ,
		x"fff821",x"fff76d",x"fff6ea",x"fff699",x"fff678",x"fff684",x"fff6ba",x"fff717" ,
		x"fff798",x"fff838",x"fff8f4",x"fff9c6",x"fffaaa",x"fffb9b",x"fffc95",x"fffd93" ,
		x"fffe91",x"ffff8a",x"00007b",x"00015f",x"000234",x"0002f5",x"0003a2",x"000437" ,
		x"0004b3",x"000515",x"00055b",x"000587",x"000598",x"00058e",x"00056c",x"000531" ,
		x"0004e1",x"00047d",x"000407",x"000383",x"0002f3",x"000259",x"0001ba",x"000118" ,
		x"000075",x"ffffd5",x"ffff3a",x"fffea8",x"fffe20",x"fffda4",x"fffd36",x"fffcd9" ,
		x"fffc8c",x"fffc52",x"fffc2a",x"fffc14",x"fffc12",x"fffc21",x"fffc42",x"fffc74" ,
		x"fffcb4",x"fffd03",x"fffd5d",x"fffdc1",x"fffe2d",x"fffe9f",x"ffff15",x"ffff8d" ,
		x"000003",x"000077",x"0000e6",x"00014f",x"0001af",x"000206",x"000251",x"000290" ,
		x"0002c1",x"0002e5",x"0002fb",x"000303",x"0002fc",x"0002e8",x"0002c7",x"000299" ,
		x"000260",x"00021e",x"0001d3",x"000181",x"00012a",x"0000cf",x"000072",x"000014" ,
		x"ffffb8",x"ffff5f",x"ffff0b",x"fffebc",x"fffe75",x"fffe36",x"fffe01",x"fffdd6" ,
		x"fffdb5",x"fffda0",x"fffd96",x"fffd98",x"fffda5",x"fffdbc",x"fffddd",x"fffe08" ,
		x"fffe3b",x"fffe76",x"fffeb7",x"fffefc",x"ffff45",x"ffff91",x"ffffdd",x"000028" ,
		x"000072",x"0000b8",x"0000fa",x"000136",x"00016c",x"00019a",x"0001c1",x"0001de" ,
		x"0001f2",x"0001fd",x"0001ff",x"0001f7",x"0001e6",x"0001cd",x"0001ac",x"000184" ,
		x"000155",x"000120",x"0000e7",x"0000ab",x"00006d",x"00002d",x"ffffee",x"ffffb0" ,
		x"ffff74",x"ffff3c",x"ffff08",x"fffed9",x"fffeb0",x"fffe8e",x"fffe73",x"fffe60" ,
		x"fffe54",x"fffe51",x"fffe55",x"fffe61",x"fffe74",x"fffe8e",x"fffeaf",x"fffed5" ,
		x"ffff00",x"ffff2f",x"ffff62",x"ffff96",x"ffffcc",x"000002",x"000037",x"00006b" ,
		x"00009b",x"0000c9",x"0000f2",x"000116",x"000135",x"00014e",x"000160",x"00016c" ,
		x"000171",x"00016f",x"000167",x"000158",x"000143",x"000129",x"000109",x"0000e6" ,
		x"0000be",x"000093",x"000067",x"000039",x"00000a",x"ffffdc",x"ffffaf",x"ffff85" ,
		x"ffff5d",x"ffff38",x"ffff17",x"fffefb",x"fffee5",x"fffed3",x"fffec7",x"fffec1" ,
		x"fffec1",x"fffec7",x"fffed2",x"fffee3",x"fffef8",x"ffff13",x"ffff31",x"ffff52" ,
		x"ffff76",x"ffff9d",x"ffffc4",x"ffffed",x"000015",x"00003c",x"000062",x"000085" ,
		x"0000a6",x"0000c3",x"0000dd",x"0000f2",x"000102",x"00010e",x"000114",x"000116" ,
		x"000112",x"00010a",x"0000fd",x"0000eb",x"0000d5",x"0000bc",x"0000a0",x"000080" ,
		x"00005f",x"00003d",x"00001a",x"fffff7",x"ffffd4",x"ffffb3",x"ffff93",x"ffff76" ,
		x"ffff5c",x"ffff44",x"ffff31",x"ffff21",x"ffff16",x"ffff0f",x"ffff0d",x"ffff0f" ,
		x"ffff15",x"ffff1f",x"ffff2e",x"ffff40",x"ffff55",x"ffff6e",x"ffff88",x"ffffa5" ,
		x"ffffc2",x"ffffe1",x"000000",x"00001e",x"00003c",x"000058",x"000073",x"00008a" ,
		x"0000a0",x"0000b2",x"0000c0",x"0000cb",x"0000d2",x"0000d6",x"0000d5",x"0000d0" ,
		x"0000c8",x"0000bc",x"0000ad",x"00009b",x"000087",x"000070",x"000057",x"00003d" ,
		x"000022",x"000007",x"ffffec",x"ffffd2",x"ffffb9",x"ffffa1",x"ffff8b",x"ffff78" ,
		x"ffff67",x"ffff5a",x"ffff4f",x"ffff48",x"ffff44",x"ffff44",x"ffff47",x"ffff4d" ,
		x"ffff57",x"ffff63",x"ffff73",x"ffff84",x"ffff98",x"ffffae",x"ffffc4",x"ffffdc" ,
		x"fffff4",x"00000c",x"000023",x"00003a",x"00004f",x"000062",x"000074",x"000083" ,
		x"000090",x"00009a",x"0000a1",x"0000a5",x"0000a7",x"0000a5",x"0000a0",x"000098" ,
		x"00008d",x"000080",x"000071",x"000060",x"00004e",x"00003a",x"000025",x"000010" ,
		x"fffffb",x"ffffe6",x"ffffd2",x"ffffbe",x"ffffad",x"ffff9d",x"ffff8e",x"ffff82" ,
		x"ffff79",x"ffff72",x"ffff6e",x"ffff6c",x"ffff6d",x"ffff71",x"ffff77",x"ffff80" ,
		x"ffff8b",x"ffff98",x"ffffa7",x"ffffb7",x"ffffc9",x"ffffdb",x"ffffee",x"000001" ,
		x"000014",x"000026",x"000037",x"000048",x"000056",x"000063",x"00006f",x"000077" ,
		x"00007e",x"000082",x"000084",x"000084",x"000081",x"00007c",x"000074",x"00006a" ,
		x"00005f",x"000052",x"000044",x"000034",x"000024",x"000012",x"000001",x"fffff1" ,
		x"ffffe0",x"ffffd0",x"ffffc1",x"ffffb4",x"ffffa7",x"ffff9c",x"ffff95",x"ffff8d" ,
		x"ffff8a",x"ffff87",x"ffff87",x"ffff8a",x"ffff8e",x"ffff95",x"ffff9e",x"ffffa8" ,
		x"ffffb4",x"ffffc1",x"ffffcf",x"ffffdf",x"ffffee",x"fffffe",x"00000e",x"00001e" ,
		x"00002d",x"00003c",x"000049",x"000054",x"00005f",x"000067",x"00006d",x"000072" ,
		x"000074",x"000074",x"000072",x"00006e",x"000068",x"000060",x"000056",x"00004a" ,
		x"00003d",x"00002e",x"00001f",x"00000f",x"ffffff",x"ffffee",x"ffffde",x"ffffce" ,
		x"ffffbf",x"ffffb1",x"ffffa4",x"ffff99",x"ffff8f",x"ffff87",x"ffff82",x"ffff7e" ,
		x"ffff7d",x"ffff7f",x"ffff82",x"ffff88",x"ffff91",x"ffff9b",x"ffffa8",x"ffffb7" ,
		x"ffffc8",x"ffffda",x"ffffee",x"000003",x"000018",x"00002f",x"000046",x"00005c" ,
		x"000073",x"000089",x"00009f",x"0000b3",x"0000c7",x"0000d8",x"0000e9",x"0000f7" ,
		x"000104",x"00010e",x"000117",x"00011d",x"000121",x"000123",x"000122",x"000120" ,
		x"00011b",x"000115",x"00010d",x"000103",x"0000f9",x"0000ed",x"0000e2",x"0000d8" ,
		x"0000d0",x"0000ce",x"0000d7",x"0000f4",x"000136",x"0001bb",x"fffe56",
		others=>x"000000"
	);
	
	constant COEFFICIENTS_6_LEN: tCoeffLenRange := 999;
	constant COEFFICIENTS_6: tCoeff := (
		x"ffffef",x"ffffec",x"ffffe9",x"ffffe7",x"ffffe5",x"ffffe3",x"ffffe2",x"ffffe2" ,
		x"ffffe2",x"ffffe2",x"ffffe3",x"ffffe5",x"ffffe7",x"ffffe9",x"ffffec",x"ffffef" ,
		x"fffff3",x"fffff7",x"fffffa",x"ffffff",x"000003",x"000007",x"00000b",x"00000f" ,
		x"000012",x"000016",x"000019",x"00001c",x"00001e",x"000020",x"000021",x"000022" ,
		x"000022",x"000021",x"000020",x"00001f",x"00001c",x"00001a",x"000016",x"000013" ,
		x"00000f",x"00000a",x"000005",x"000001",x"fffffc",x"fffff7",x"fffff2",x"ffffed" ,
		x"ffffe8",x"ffffe4",x"ffffe0",x"ffffdc",x"ffffda",x"ffffd7",x"ffffd6",x"ffffd5" ,
		x"ffffd4",x"ffffd5",x"ffffd6",x"ffffd8",x"ffffdb",x"ffffde",x"ffffe2",x"ffffe7" ,
		x"ffffec",x"fffff2",x"fffff8",x"fffffe",x"000005",x"00000b",x"000012",x"000018" ,
		x"00001e",x"000024",x"000029",x"00002d",x"000031",x"000034",x"000037",x"000038" ,
		x"000038",x"000038",x"000036",x"000034",x"000030",x"00002c",x"000026",x"000020" ,
		x"000019",x"000012",x"00000a",x"000001",x"fffff9",x"fffff0",x"ffffe7",x"ffffdf" ,
		x"ffffd7",x"ffffcf",x"ffffc8",x"ffffc2",x"ffffbd",x"ffffb9",x"ffffb6",x"ffffb4" ,
		x"ffffb3",x"ffffb4",x"ffffb6",x"ffffba",x"ffffbe",x"ffffc4",x"ffffcc",x"ffffd4" ,
		x"ffffdd",x"ffffe7",x"fffff2",x"fffffd",x"000009",x"000015",x"000020",x"00002c" ,
		x"000036",x"000040",x"00004a",x"000052",x"000059",x"00005e",x"000062",x"000065" ,
		x"000065",x"000064",x"000061",x"00005d",x"000056",x"00004e",x"000044",x"000039" ,
		x"00002d",x"00001f",x"000011",x"000002",x"fffff3",x"ffffe3",x"ffffd4",x"ffffc5" ,
		x"ffffb7",x"ffffa9",x"ffff9d",x"ffff92",x"ffff89",x"ffff82",x"ffff7d",x"ffff7a" ,
		x"ffff79",x"ffff7b",x"ffff7f",x"ffff85",x"ffff8e",x"ffff98",x"ffffa5",x"ffffb4" ,
		x"ffffc4",x"ffffd6",x"ffffe9",x"fffffc",x"000010",x"000025",x"000039",x"00004c" ,
		x"00005f",x"000070",x"000080",x"00008e",x"00009a",x"0000a3",x"0000a9",x"0000ad" ,
		x"0000ae",x"0000ac",x"0000a7",x"00009e",x"000093",x"000085",x"000074",x"000061" ,
		x"00004c",x"000035",x"00001d",x"000003",x"ffffe9",x"ffffcf",x"ffffb5",x"ffff9c" ,
		x"ffff84",x"ffff6e",x"ffff5a",x"ffff48",x"ffff39",x"ffff2e",x"ffff25",x"ffff20" ,
		x"ffff20",x"ffff23",x"ffff29",x"ffff34",x"ffff43",x"ffff55",x"ffff6a",x"ffff83" ,
		x"ffff9e",x"ffffbb",x"ffffda",x"fffffb",x"00001c",x"00003d",x"00005e",x"00007e" ,
		x"00009d",x"0000b9",x"0000d2",x"0000e9",x"0000fb",x"00010a",x"000115",x"00011a" ,
		x"00011b",x"000117",x"00010e",x"000101",x"0000ee",x"0000d7",x"0000bc",x"00009d" ,
		x"00007a",x"000055",x"00002e",x"000005",x"ffffdb",x"ffffb1",x"ffff88",x"ffff5f" ,
		x"ffff39",x"ffff16",x"fffef6",x"fffeda",x"fffec3",x"fffeb0",x"fffea3",x"fffe9c" ,
		x"fffe9b",x"fffea0",x"fffeac",x"fffebd",x"fffed5",x"fffef2",x"ffff14",x"ffff3b" ,
		x"ffff66",x"ffff95",x"ffffc6",x"fffff9",x"00002e",x"000062",x"000096",x"0000c8" ,
		x"0000f8",x"000124",x"00014b",x"00016e",x"00018b",x"0001a2",x"0001b2",x"0001ba" ,
		x"0001bc",x"0001b5",x"0001a7",x"000191",x"000173",x"00014f",x"000124",x"0000f3" ,
		x"0000be",x"000084",x"000046",x"000006",x"ffffc5",x"ffff84",x"ffff44",x"ffff06" ,
		x"fffecb",x"fffe94",x"fffe62",x"fffe37",x"fffe13",x"fffdf7",x"fffde4",x"fffdd9" ,
		x"fffdd8",x"fffde1",x"fffdf2",x"fffe0e",x"fffe32",x"fffe60",x"fffe95",x"fffed1" ,
		x"ffff14",x"ffff5c",x"ffffa9",x"fffff8",x"000049",x"00009a",x"0000e9",x"000137" ,
		x"000180",x"0001c4",x"000201",x"000236",x"000263",x"000286",x"00029e",x"0002ab" ,
		x"0002ac",x"0002a2",x"00028b",x"000269",x"00023c",x"000204",x"0001c1",x"000176" ,
		x"000123",x"0000c9",x"00006a",x"000008",x"ffffa3",x"ffff3e",x"fffedb",x"fffe7b" ,
		x"fffe20",x"fffdcb",x"fffd7f",x"fffd3c",x"fffd05",x"fffcd9",x"fffcbb",x"fffcab" ,
		x"fffca9",x"fffcb6",x"fffcd2",x"fffcfc",x"fffd35",x"fffd7b",x"fffdce",x"fffe2c" ,
		x"fffe94",x"ffff04",x"ffff7b",x"fffff7",x"000075",x"0000f3",x"000170",x"0001e9" ,
		x"00025c",x"0002c6",x"000326",x"00037b",x"0003c1",x"0003f8",x"00041f",x"000434" ,
		x"000437",x"000427",x"000404",x"0003cf",x"000387",x"00032f",x"0002c7",x"000250" ,
		x"0001cc",x"00013d",x"0000a6",x"000009",x"ffff68",x"fffec7",x"fffe27",x"fffd8c" ,
		x"fffcf9",x"fffc70",x"fffbf3",x"fffb86",x"fffb2b",x"fffae3",x"fffab0",x"fffa93" ,
		x"fffa8e",x"fffaa1",x"fffacd",x"fffb10",x"fffb6b",x"fffbdd",x"fffc64",x"fffcfe" ,
		x"fffda9",x"fffe62",x"ffff28",x"fffff6",x"0000c9",x"00019e",x"000271",x"00033e" ,
		x"000403",x"0004ba",x"000561",x"0005f5",x"000672",x"0006d5",x"00071d",x"000746" ,
		x"000751",x"00073b",x"000704",x"0006ad",x"000635",x"00059e",x"0004ea",x"00041a" ,
		x"000332",x"000235",x"000126",x"00000a",x"fffee5",x"fffdbb",x"fffc93",x"fffb70" ,
		x"fffa58",x"fff950",x"fff85e",x"fff785",x"fff6cb",x"fff633",x"fff5c3",x"fff57c" ,
		x"fff561",x"fff575",x"fff5b9",x"fff62e",x"fff6d3",x"fff7a8",x"fff8ab",x"fff9d9" ,
		x"fffb2f",x"fffca9",x"fffe42",x"fffff5",x"0001bb",x"00038f",x"000567",x"00073e" ,
		x"00090b",x"000ac5",x"000c66",x"000de3",x"000f37",x"001058",x"00113f",x"0011e5" ,
		x"001244",x"001256",x"001216",x"001180",x"001090",x"000f45",x"000d9d",x"000b98" ,
		x"000937",x"00067d",x"00036c",x"00000a",x"fffc5b",x"fff867",x"fff434",x"ffefcc" ,
		x"ffeb36",x"ffe67e",x"ffe1ae",x"ffdcd1",x"ffd7f2",x"ffd31c",x"ffce5d",x"ffc9be" ,
		x"ffc54d",x"ffc113",x"ffbd1d",x"ffb973",x"ffb61f",x"ffb32b",x"ffb09d",x"ffae7d" ,
		x"ffaccf",x"ffab99",x"ffaade",x"07aaa0",x"ffaade",x"ffab99",x"ffaccf",x"ffae7d" ,
		x"ffb09d",x"ffb32b",x"ffb61f",x"ffb973",x"ffbd1d",x"ffc113",x"ffc54d",x"ffc9be" ,
		x"ffce5d",x"ffd31c",x"ffd7f2",x"ffdcd1",x"ffe1ae",x"ffe67e",x"ffeb36",x"ffefcc" ,
		x"fff434",x"fff867",x"fffc5b",x"00000a",x"00036c",x"00067d",x"000937",x"000b98" ,
		x"000d9d",x"000f45",x"001090",x"001180",x"001216",x"001256",x"001244",x"0011e5" ,
		x"00113f",x"001058",x"000f37",x"000de3",x"000c66",x"000ac5",x"00090b",x"00073e" ,
		x"000567",x"00038f",x"0001bb",x"fffff5",x"fffe42",x"fffca9",x"fffb2f",x"fff9d9" ,
		x"fff8ab",x"fff7a8",x"fff6d3",x"fff62e",x"fff5b9",x"fff575",x"fff561",x"fff57c" ,
		x"fff5c3",x"fff633",x"fff6cb",x"fff785",x"fff85e",x"fff950",x"fffa58",x"fffb70" ,
		x"fffc93",x"fffdbb",x"fffee5",x"00000a",x"000126",x"000235",x"000332",x"00041a" ,
		x"0004ea",x"00059e",x"000635",x"0006ad",x"000704",x"00073b",x"000751",x"000746" ,
		x"00071d",x"0006d5",x"000672",x"0005f5",x"000561",x"0004ba",x"000403",x"00033e" ,
		x"000271",x"00019e",x"0000c9",x"fffff6",x"ffff28",x"fffe62",x"fffda9",x"fffcfe" ,
		x"fffc64",x"fffbdd",x"fffb6b",x"fffb10",x"fffacd",x"fffaa1",x"fffa8e",x"fffa93" ,
		x"fffab0",x"fffae3",x"fffb2b",x"fffb86",x"fffbf3",x"fffc70",x"fffcf9",x"fffd8c" ,
		x"fffe27",x"fffec7",x"ffff68",x"000009",x"0000a6",x"00013d",x"0001cc",x"000250" ,
		x"0002c7",x"00032f",x"000387",x"0003cf",x"000404",x"000427",x"000437",x"000434" ,
		x"00041f",x"0003f8",x"0003c1",x"00037b",x"000326",x"0002c6",x"00025c",x"0001e9" ,
		x"000170",x"0000f3",x"000075",x"fffff7",x"ffff7b",x"ffff04",x"fffe94",x"fffe2c" ,
		x"fffdce",x"fffd7b",x"fffd35",x"fffcfc",x"fffcd2",x"fffcb6",x"fffca9",x"fffcab" ,
		x"fffcbb",x"fffcd9",x"fffd05",x"fffd3c",x"fffd7f",x"fffdcb",x"fffe20",x"fffe7b" ,
		x"fffedb",x"ffff3e",x"ffffa3",x"000008",x"00006a",x"0000c9",x"000123",x"000176" ,
		x"0001c1",x"000204",x"00023c",x"000269",x"00028b",x"0002a2",x"0002ac",x"0002ab" ,
		x"00029e",x"000286",x"000263",x"000236",x"000201",x"0001c4",x"000180",x"000137" ,
		x"0000e9",x"00009a",x"000049",x"fffff8",x"ffffa9",x"ffff5c",x"ffff14",x"fffed1" ,
		x"fffe95",x"fffe60",x"fffe32",x"fffe0e",x"fffdf2",x"fffde1",x"fffdd8",x"fffdd9" ,
		x"fffde4",x"fffdf7",x"fffe13",x"fffe37",x"fffe62",x"fffe94",x"fffecb",x"ffff06" ,
		x"ffff44",x"ffff84",x"ffffc5",x"000006",x"000046",x"000084",x"0000be",x"0000f3" ,
		x"000124",x"00014f",x"000173",x"000191",x"0001a7",x"0001b5",x"0001bc",x"0001ba" ,
		x"0001b2",x"0001a2",x"00018b",x"00016e",x"00014b",x"000124",x"0000f8",x"0000c8" ,
		x"000096",x"000062",x"00002e",x"fffff9",x"ffffc6",x"ffff95",x"ffff66",x"ffff3b" ,
		x"ffff14",x"fffef2",x"fffed5",x"fffebd",x"fffeac",x"fffea0",x"fffe9b",x"fffe9c" ,
		x"fffea3",x"fffeb0",x"fffec3",x"fffeda",x"fffef6",x"ffff16",x"ffff39",x"ffff5f" ,
		x"ffff88",x"ffffb1",x"ffffdb",x"000005",x"00002e",x"000055",x"00007a",x"00009d" ,
		x"0000bc",x"0000d7",x"0000ee",x"000101",x"00010e",x"000117",x"00011b",x"00011a" ,
		x"000115",x"00010a",x"0000fb",x"0000e9",x"0000d2",x"0000b9",x"00009d",x"00007e" ,
		x"00005e",x"00003d",x"00001c",x"fffffb",x"ffffda",x"ffffbb",x"ffff9e",x"ffff83" ,
		x"ffff6a",x"ffff55",x"ffff43",x"ffff34",x"ffff29",x"ffff23",x"ffff20",x"ffff20" ,
		x"ffff25",x"ffff2e",x"ffff39",x"ffff48",x"ffff5a",x"ffff6e",x"ffff84",x"ffff9c" ,
		x"ffffb5",x"ffffcf",x"ffffe9",x"000003",x"00001d",x"000035",x"00004c",x"000061" ,
		x"000074",x"000085",x"000093",x"00009e",x"0000a7",x"0000ac",x"0000ae",x"0000ad" ,
		x"0000a9",x"0000a3",x"00009a",x"00008e",x"000080",x"000070",x"00005f",x"00004c" ,
		x"000039",x"000025",x"000010",x"fffffc",x"ffffe9",x"ffffd6",x"ffffc4",x"ffffb4" ,
		x"ffffa5",x"ffff98",x"ffff8e",x"ffff85",x"ffff7f",x"ffff7b",x"ffff79",x"ffff7a" ,
		x"ffff7d",x"ffff82",x"ffff89",x"ffff92",x"ffff9d",x"ffffa9",x"ffffb7",x"ffffc5" ,
		x"ffffd4",x"ffffe3",x"fffff3",x"000002",x"000011",x"00001f",x"00002d",x"000039" ,
		x"000044",x"00004e",x"000056",x"00005d",x"000061",x"000064",x"000065",x"000065" ,
		x"000062",x"00005e",x"000059",x"000052",x"00004a",x"000040",x"000036",x"00002c" ,
		x"000020",x"000015",x"000009",x"fffffd",x"fffff2",x"ffffe7",x"ffffdd",x"ffffd4" ,
		x"ffffcc",x"ffffc4",x"ffffbe",x"ffffba",x"ffffb6",x"ffffb4",x"ffffb3",x"ffffb4" ,
		x"ffffb6",x"ffffb9",x"ffffbd",x"ffffc2",x"ffffc8",x"ffffcf",x"ffffd7",x"ffffdf" ,
		x"ffffe7",x"fffff0",x"fffff9",x"000001",x"00000a",x"000012",x"000019",x"000020" ,
		x"000026",x"00002c",x"000030",x"000034",x"000036",x"000038",x"000038",x"000038" ,
		x"000037",x"000034",x"000031",x"00002d",x"000029",x"000024",x"00001e",x"000018" ,
		x"000012",x"00000b",x"000005",x"fffffe",x"fffff8",x"fffff2",x"ffffec",x"ffffe7" ,
		x"ffffe2",x"ffffde",x"ffffdb",x"ffffd8",x"ffffd6",x"ffffd5",x"ffffd4",x"ffffd5" ,
		x"ffffd6",x"ffffd7",x"ffffda",x"ffffdc",x"ffffe0",x"ffffe4",x"ffffe8",x"ffffed" ,
		x"fffff2",x"fffff7",x"fffffc",x"000001",x"000005",x"00000a",x"00000f",x"000013" ,
		x"000016",x"00001a",x"00001c",x"00001f",x"000020",x"000021",x"000022",x"000022" ,
		x"000021",x"000020",x"00001e",x"00001c",x"000019",x"000016",x"000012",x"00000f" ,
		x"00000b",x"000007",x"000003",x"ffffff",x"fffffa",x"fffff7",x"fffff3",x"ffffef" ,
		x"ffffec",x"ffffe9",x"ffffe7",x"ffffe5",x"ffffe3",x"ffffe2",x"ffffe2",x"ffffe2" ,
		x"ffffe2",x"ffffe3",x"ffffe5",x"ffffe7",x"ffffe9",x"ffffec",x"ffffef",
		others=>x"000000"
	);
	
	constant COEFFICIENTS_7_LEN: tCoeffLenRange := 999;
	constant COEFFICIENTS_7: tCoeff := (
		x"ffffd2",x"ffffce",x"ffffcd",x"ffffce",x"ffffd1",x"ffffd5",x"ffffdc",x"ffffe3" ,
		x"ffffea",x"fffff2",x"fffff9",x"000000",x"000004",x"000008",x"000009",x"000009" ,
		x"000008",x"000005",x"000002",x"fffffe",x"fffffa",x"fffff6",x"fffff4",x"fffff2" ,
		x"fffff3",x"fffff5",x"fffff9",x"ffffff",x"000007",x"000010",x"000019",x"000023" ,
		x"00002c",x"000034",x"00003a",x"00003e",x"00003f",x"00003e",x"000039",x"000032" ,
		x"000028",x"00001c",x"00000e",x"000000",x"fffff1",x"ffffe2",x"ffffd5",x"ffffca" ,
		x"ffffc1",x"ffffbc",x"ffffb9",x"ffffb9",x"ffffbd",x"ffffc3",x"ffffcc",x"ffffd6" ,
		x"ffffe1",x"ffffec",x"fffff6",x"ffffff",x"000007",x"00000c",x"00000f",x"00000f" ,
		x"00000d",x"000009",x"000003",x"fffffd",x"fffff6",x"fffff1",x"ffffed",x"ffffeb" ,
		x"ffffeb",x"ffffef",x"fffff6",x"000000",x"00000c",x"00001a",x"00002a",x"00003a" ,
		x"000049",x"000056",x"000061",x"000068",x"00006b",x"000068",x"000061",x"000055" ,
		x"000045",x"000030",x"000019",x"000000",x"ffffe6",x"ffffcd",x"ffffb6",x"ffffa2" ,
		x"ffff93",x"ffff89",x"ffff84",x"ffff84",x"ffff8a",x"ffff95",x"ffffa4",x"ffffb6" ,
		x"ffffc9",x"ffffdd",x"ffffef",x"ffffff",x"00000d",x"000016",x"00001b",x"00001b" ,
		x"000018",x"000010",x"000006",x"fffffb",x"fffff0",x"ffffe6",x"ffffde",x"ffffdb" ,
		x"ffffdc",x"ffffe2",x"ffffee",x"000000",x"000015",x"00002f",x"00004b",x"000067" ,
		x"000082",x"00009a",x"0000ad",x"0000ba",x"0000be",x"0000bb",x"0000ae",x"000098" ,
		x"00007b",x"000056",x"00002c",x"ffffff",x"ffffd2",x"ffffa5",x"ffff7d",x"ffff5a" ,
		x"ffff3f",x"ffff2d",x"ffff24",x"ffff25",x"ffff30",x"ffff44",x"ffff5e",x"ffff7d" ,
		x"ffff9f",x"ffffc2",x"ffffe3",x"000000",x"000017",x"000027",x"000030",x"000031" ,
		x"00002a",x"00001e",x"00000c",x"fffff9",x"ffffe5",x"ffffd4",x"ffffc7",x"ffffc1" ,
		x"ffffc2",x"ffffcd",x"ffffe2",x"ffffff",x"000025",x"000051",x"000080",x"0000b1" ,
		x"0000df",x"000108",x"000128",x"00013d",x"000145",x"00013e",x"000128",x"000103" ,
		x"0000d1",x"000092",x"00004c",x"000000",x"ffffb2",x"ffff67",x"ffff23",x"fffee8" ,
		x"fffebb",x"fffe9c",x"fffe8e",x"fffe91",x"fffea3",x"fffec4",x"fffef0",x"ffff25" ,
		x"ffff5e",x"ffff98",x"ffffcf",x"ffffff",x"000026",x"000042",x"000050",x"000052" ,
		x"000047",x"000033",x"000016",x"fffff6",x"ffffd6",x"ffffb9",x"ffffa4",x"ffff99" ,
		x"ffff9c",x"ffffae",x"ffffcf",x"000000",x"00003d",x"000084",x"0000d1",x"00011f" ,
		x"00016a",x"0001ac",x"0001e0",x"000202",x"00020e",x"000203",x"0001df",x"0001a3" ,
		x"000151",x"0000ec",x"00007a",x"ffffff",x"ffff83",x"ffff0b",x"fffe9d",x"fffe3f" ,
		x"fffdf7",x"fffdc6",x"fffdb0",x"fffdb4",x"fffdd2",x"fffe07",x"fffe4e",x"fffea2" ,
		x"fffefe",x"ffff5a",x"ffffb2",x"000000",x"00003e",x"000069",x"000081",x"000083" ,
		x"000073",x"000052",x"000026",x"fffff3",x"ffffc0",x"ffff93",x"ffff71",x"ffff60" ,
		x"ffff64",x"ffff80",x"ffffb4",x"000000",x"00005f",x"0000ce",x"000146",x"0001c1" ,
		x"000236",x"00029c",x"0002ed",x"000322",x"000335",x"000323",x"0002ea",x"00028d" ,
		x"00020d",x"000170",x"0000be",x"ffffff",x"ffff3e",x"fffe83",x"fffdd8",x"fffd47" ,
		x"fffcd6",x"fffc8b",x"fffc68",x"fffc6f",x"fffc9e",x"fffcef",x"fffd5e",x"fffde0" ,
		x"fffe6f",x"fffeff",x"ffff87",x"000000",x"000060",x"0000a4",x"0000c9",x"0000ce" ,
		x"0000b5",x"000083",x"00003f",x"fffff0",x"ffffa1",x"ffff5b",x"ffff27",x"ffff0c" ,
		x"ffff12",x"ffff3d",x"ffff8c",x"ffffff",x"000092",x"00013d",x"0001f6",x"0002b3" ,
		x"000366",x"000404",x"000481",x"0004d3",x"0004f1",x"0004d5",x"00047f",x"0003ef" ,
		x"00032a",x"000238",x"000126",x"000000",x"fffed4",x"fffdb3",x"fffcab",x"fffbca" ,
		x"fffb1a",x"fffaa5",x"fffa6f",x"fffa79",x"fffac1",x"fffb3e",x"fffbe9",x"fffcb3" ,
		x"fffd90",x"fffe70",x"ffff44",x"ffffff",x"000097",x"000102",x"00013c",x"000144" ,
		x"00011f",x"0000d2",x"000068",x"ffffee",x"ffff72",x"ffff04",x"fffeb2",x"fffe87" ,
		x"fffe90",x"fffed0",x"ffff4c",x"000000",x"0000e5",x"0001f0",x"000314",x"00043d" ,
		x"000559",x"000654",x"00071b",x"00079e",x"0007d0",x"0007a7",x"000721",x"00063e" ,
		x"000508",x"000389",x"0001d5",x"ffffff",x"fffe20",x"fffc50",x"fffaa7",x"fff93a" ,
		x"fff81d",x"fff75c",x"fff701",x"fff70d",x"fff77c",x"fff844",x"fff955",x"fffa9d" ,
		x"fffc03",x"fffd70",x"fffecb",x"000000",x"0000fa",x"0001ac",x"00020f",x"000220" ,
		x"0001e4",x"000166",x"0000b7",x"ffffec",x"ffff1d",x"fffe63",x"fffdd6",x"fffd8b" ,
		x"fffd96",x"fffe00",x"fffecf",x"ffffff",x"000187",x"000353",x"00054a",x"000750" ,
		x"000943",x"000b01",x"000c68",x"000d5a",x"000dbf",x"000d86",x"000ca6",x"000b21" ,
		x"000902",x"00065d",x"000350",x"000000",x"fffc96",x"fff93e",x"fff626",x"fff375" ,
		x"fff150",x"ffefd2",x"ffef0e",x"ffef0a",x"ffefc3",x"fff129",x"fff320",x"fff586" ,
		x"fff830",x"fffaf1",x"fffd9b",x"ffffff",x"0001f9",x"00036a",x"00043d",x"00046c" ,
		x"0003fb",x"0002ff",x"000197",x"ffffeb",x"fffe2d",x"fffc92",x"fffb51",x"fffa9d" ,
		x"fffaa1",x"fffb7f",x"fffd48",x"000000",x"000396",x"0007ea",x"000cc8",x"0011f0" ,
		x"001713",x"001bdc",x"001ff2",x"002300",x"0024b6",x"0024d2",x"002326",x"001f98" ,
		x"001a25",x"0012e9",x"000a18",x"ffffff",x"fff504",x"ffe99e",x"ffde50",x"ffd3a6" ,
		x"ffca2b",x"ffc262",x"ffbcbf",x"ffb9a2",x"ffb94e",x"ffbbe8",x"ffc172",x"ffc9c9" ,
		x"ffd4aa",x"ffe1ad",x"fff052",x"ffffff",x"00100c",x"001fc8",x"002e83",x"003b96" ,
		x"00466c",x"004e88",x"00538d",x"005540",x"00538d",x"004e88",x"00466c",x"003b96" ,
		x"002e83",x"001fc8",x"00100c",x"ffffff",x"fff052",x"ffe1ad",x"ffd4aa",x"ffc9c9" ,
		x"ffc172",x"ffbbe8",x"ffb94e",x"ffb9a2",x"ffbcbf",x"ffc262",x"ffca2b",x"ffd3a6" ,
		x"ffde50",x"ffe99e",x"fff504",x"ffffff",x"000a18",x"0012e9",x"001a25",x"001f98" ,
		x"002326",x"0024d2",x"0024b6",x"002300",x"001ff2",x"001bdc",x"001713",x"0011f0" ,
		x"000cc8",x"0007ea",x"000396",x"000000",x"fffd48",x"fffb7f",x"fffaa1",x"fffa9d" ,
		x"fffb51",x"fffc92",x"fffe2d",x"ffffeb",x"000197",x"0002ff",x"0003fb",x"00046c" ,
		x"00043d",x"00036a",x"0001f9",x"ffffff",x"fffd9b",x"fffaf1",x"fff830",x"fff586" ,
		x"fff320",x"fff129",x"ffefc3",x"ffef0a",x"ffef0e",x"ffefd2",x"fff150",x"fff375" ,
		x"fff626",x"fff93e",x"fffc96",x"000000",x"000350",x"00065d",x"000902",x"000b21" ,
		x"000ca6",x"000d86",x"000dbf",x"000d5a",x"000c68",x"000b01",x"000943",x"000750" ,
		x"00054a",x"000353",x"000187",x"ffffff",x"fffecf",x"fffe00",x"fffd96",x"fffd8b" ,
		x"fffdd6",x"fffe63",x"ffff1d",x"ffffec",x"0000b7",x"000166",x"0001e4",x"000220" ,
		x"00020f",x"0001ac",x"0000fa",x"000000",x"fffecb",x"fffd70",x"fffc03",x"fffa9d" ,
		x"fff955",x"fff844",x"fff77c",x"fff70d",x"fff701",x"fff75c",x"fff81d",x"fff93a" ,
		x"fffaa7",x"fffc50",x"fffe20",x"ffffff",x"0001d5",x"000389",x"000508",x"00063e" ,
		x"000721",x"0007a7",x"0007d0",x"00079e",x"00071b",x"000654",x"000559",x"00043d" ,
		x"000314",x"0001f0",x"0000e5",x"000000",x"ffff4c",x"fffed0",x"fffe90",x"fffe87" ,
		x"fffeb2",x"ffff04",x"ffff72",x"ffffee",x"000068",x"0000d2",x"00011f",x"000144" ,
		x"00013c",x"000102",x"000097",x"ffffff",x"ffff44",x"fffe70",x"fffd90",x"fffcb3" ,
		x"fffbe9",x"fffb3e",x"fffac1",x"fffa79",x"fffa6f",x"fffaa5",x"fffb1a",x"fffbca" ,
		x"fffcab",x"fffdb3",x"fffed4",x"000000",x"000126",x"000238",x"00032a",x"0003ef" ,
		x"00047f",x"0004d5",x"0004f1",x"0004d3",x"000481",x"000404",x"000366",x"0002b3" ,
		x"0001f6",x"00013d",x"000092",x"ffffff",x"ffff8c",x"ffff3d",x"ffff12",x"ffff0c" ,
		x"ffff27",x"ffff5b",x"ffffa1",x"fffff0",x"00003f",x"000083",x"0000b5",x"0000ce" ,
		x"0000c9",x"0000a4",x"000060",x"000000",x"ffff87",x"fffeff",x"fffe6f",x"fffde0" ,
		x"fffd5e",x"fffcef",x"fffc9e",x"fffc6f",x"fffc68",x"fffc8b",x"fffcd6",x"fffd47" ,
		x"fffdd8",x"fffe83",x"ffff3e",x"ffffff",x"0000be",x"000170",x"00020d",x"00028d" ,
		x"0002ea",x"000323",x"000335",x"000322",x"0002ed",x"00029c",x"000236",x"0001c1" ,
		x"000146",x"0000ce",x"00005f",x"000000",x"ffffb4",x"ffff80",x"ffff64",x"ffff60" ,
		x"ffff71",x"ffff93",x"ffffc0",x"fffff3",x"000026",x"000052",x"000073",x"000083" ,
		x"000081",x"000069",x"00003e",x"000000",x"ffffb2",x"ffff5a",x"fffefe",x"fffea2" ,
		x"fffe4e",x"fffe07",x"fffdd2",x"fffdb4",x"fffdb0",x"fffdc6",x"fffdf7",x"fffe3f" ,
		x"fffe9d",x"ffff0b",x"ffff83",x"ffffff",x"00007a",x"0000ec",x"000151",x"0001a3" ,
		x"0001df",x"000203",x"00020e",x"000202",x"0001e0",x"0001ac",x"00016a",x"00011f" ,
		x"0000d1",x"000084",x"00003d",x"000000",x"ffffcf",x"ffffae",x"ffff9c",x"ffff99" ,
		x"ffffa4",x"ffffb9",x"ffffd6",x"fffff6",x"000016",x"000033",x"000047",x"000052" ,
		x"000050",x"000042",x"000026",x"ffffff",x"ffffcf",x"ffff98",x"ffff5e",x"ffff25" ,
		x"fffef0",x"fffec4",x"fffea3",x"fffe91",x"fffe8e",x"fffe9c",x"fffebb",x"fffee8" ,
		x"ffff23",x"ffff67",x"ffffb2",x"000000",x"00004c",x"000092",x"0000d1",x"000103" ,
		x"000128",x"00013e",x"000145",x"00013d",x"000128",x"000108",x"0000df",x"0000b1" ,
		x"000080",x"000051",x"000025",x"ffffff",x"ffffe2",x"ffffcd",x"ffffc2",x"ffffc1" ,
		x"ffffc7",x"ffffd4",x"ffffe5",x"fffff9",x"00000c",x"00001e",x"00002a",x"000031" ,
		x"000030",x"000027",x"000017",x"000000",x"ffffe3",x"ffffc2",x"ffff9f",x"ffff7d" ,
		x"ffff5e",x"ffff44",x"ffff30",x"ffff25",x"ffff24",x"ffff2d",x"ffff3f",x"ffff5a" ,
		x"ffff7d",x"ffffa5",x"ffffd2",x"ffffff",x"00002c",x"000056",x"00007b",x"000098" ,
		x"0000ae",x"0000bb",x"0000be",x"0000ba",x"0000ad",x"00009a",x"000082",x"000067" ,
		x"00004b",x"00002f",x"000015",x"000000",x"ffffee",x"ffffe2",x"ffffdc",x"ffffdb" ,
		x"ffffde",x"ffffe6",x"fffff0",x"fffffb",x"000006",x"000010",x"000018",x"00001b" ,
		x"00001b",x"000016",x"00000d",x"ffffff",x"ffffef",x"ffffdd",x"ffffc9",x"ffffb6" ,
		x"ffffa4",x"ffff95",x"ffff8a",x"ffff84",x"ffff84",x"ffff89",x"ffff93",x"ffffa2" ,
		x"ffffb6",x"ffffcd",x"ffffe6",x"000000",x"000019",x"000030",x"000045",x"000055" ,
		x"000061",x"000068",x"00006b",x"000068",x"000061",x"000056",x"000049",x"00003a" ,
		x"00002a",x"00001a",x"00000c",x"000000",x"fffff6",x"ffffef",x"ffffeb",x"ffffeb" ,
		x"ffffed",x"fffff1",x"fffff6",x"fffffd",x"000003",x"000009",x"00000d",x"00000f" ,
		x"00000f",x"00000c",x"000007",x"ffffff",x"fffff6",x"ffffec",x"ffffe1",x"ffffd6" ,
		x"ffffcc",x"ffffc3",x"ffffbd",x"ffffb9",x"ffffb9",x"ffffbc",x"ffffc1",x"ffffca" ,
		x"ffffd5",x"ffffe2",x"fffff1",x"000000",x"00000e",x"00001c",x"000028",x"000032" ,
		x"000039",x"00003e",x"00003f",x"00003e",x"00003a",x"000034",x"00002c",x"000023" ,
		x"000019",x"000010",x"000007",x"ffffff",x"fffff9",x"fffff5",x"fffff3",x"fffff2" ,
		x"fffff4",x"fffff6",x"fffffa",x"fffffe",x"000002",x"000005",x"000008",x"000009" ,
		x"000009",x"000008",x"000004",x"000000",x"fffff9",x"fffff2",x"ffffea",x"ffffe3" ,
		x"ffffdc",x"ffffd5",x"ffffd1",x"ffffce",x"ffffcd",x"ffffce",x"ffffd2",
		others=>x"000000"	
	);
	
	
	
	
	
	
	
	
	
	
	constant COEFFICIENTS_8_LEN: tCoeffLenRange := 999;
	constant COEFFICIENTS_8: tCoeff := (
	x"000023",x"000021",x"00001f",x"00001b",x"000017",x"000013",x"00000f",x"00000a" ,
x"000006",x"000002",x"ffffff",x"fffffc",x"fffffa",x"fffff8",x"fffff8",x"fffff8" ,
x"fffff9",x"fffffa",x"fffffb",x"fffffd",x"ffffff",x"000001",x"000003",x"000005" ,
x"000006",x"000006",x"000005",x"000004",x"000002",x"ffffff",x"fffffc",x"fffff8" ,
x"fffff3",x"ffffee",x"ffffe9",x"ffffe4",x"ffffdf",x"ffffdb",x"ffffd7",x"ffffd5" ,
x"ffffd4",x"ffffd4",x"ffffd6",x"ffffd9",x"ffffde",x"ffffe4",x"ffffeb",x"fffff4" ,
x"fffffe",x"000009",x"000014",x"00001f",x"00002a",x"000035",x"00003e",x"000046" ,
x"00004d",x"000051",x"000053",x"000053",x"000051",x"00004c",x"000045",x"00003c" ,
x"000030",x"000023",x"000014",x"000004",x"fffff4",x"ffffe4",x"ffffd4",x"ffffc5" ,
x"ffffb8",x"ffffac",x"ffffa3",x"ffff9c",x"ffff97",x"ffff96",x"ffff97",x"ffff9c" ,
x"ffffa3",x"ffffad",x"ffffb9",x"ffffc7",x"ffffd6",x"ffffe7",x"fffff7",x"000008" ,
x"000018",x"000027",x"000034",x"000040",x"000049",x"00004f",x"000053",x"000055" ,
x"000054",x"000050",x"00004a",x"000043",x"00003a",x"00002f",x"000025",x"00001a" ,
x"00000f",x"000005",x"fffffd",x"fffff6",x"fffff0",x"ffffed",x"ffffeb",x"ffffeb" ,
x"ffffed",x"fffff1",x"fffff5",x"fffffb",x"000000",x"000006",x"00000b",x"00000f" ,
x"000012",x"000012",x"000011",x"00000d",x"000007",x"fffffe",x"fffff3",x"ffffe7" ,
x"ffffd8",x"ffffc9",x"ffffba",x"ffffaa",x"ffff9c",x"ffff8f",x"ffff85",x"ffff7d" ,
x"ffff7a",x"ffff7a",x"ffff80",x"ffff8a",x"ffff98",x"ffffac",x"ffffc3",x"ffffdf" ,
x"fffffe",x"00001f",x"000042",x"000065",x"000087",x"0000a7",x"0000c4",x"0000dd" ,
x"0000f1",x"0000fe",x"000105",x"000105",x"0000fd",x"0000ed",x"0000d6",x"0000b8" ,
x"000094",x"00006a",x"00003c",x"00000b",x"ffffd9",x"ffffa7",x"ffff76",x"ffff48" ,
x"ffff1f",x"fffefc",x"fffedf",x"fffeca",x"fffebe",x"fffebb",x"fffec1",x"fffed0" ,
x"fffee7",x"ffff06",x"ffff2b",x"ffff57",x"ffff86",x"ffffb8",x"ffffea",x"00001c" ,
x"00004d",x"000079",x"0000a0",x"0000c2",x"0000dc",x"0000ef",x"0000fa",x"0000fd" ,
x"0000f9",x"0000ed",x"0000db",x"0000c4",x"0000a8",x"00008a",x"00006a",x"00004a" ,
x"00002b",x"00000f",x"fffff6",x"ffffe2",x"ffffd3",x"ffffc9",x"ffffc5",x"ffffc7" ,
x"ffffcd",x"ffffd7",x"ffffe5",x"fffff5",x"000005",x"000015",x"000023",x"00002e" ,
x"000035",x"000036",x"000031",x"000025",x"000013",x"fffffa",x"ffffdb",x"ffffb7" ,
x"ffff8f",x"ffff64",x"ffff39",x"ffff0e",x"fffee7",x"fffec5",x"fffeaa",x"fffe97" ,
x"fffe8f",x"fffe93",x"fffea3",x"fffebf",x"fffee9",x"ffff20",x"ffff62",x"ffffae" ,
x"000002",x"00005b",x"0000b9",x"000116",x"000171",x"0001c5",x"000211",x"000252" ,
x"000284",x"0002a5",x"0002b5",x"0002b1",x"000298",x"00026c",x"00022d",x"0001dc" ,
x"00017b",x"00010d",x"000094",x"000014",x"ffff92",x"ffff10",x"fffe93",x"fffe1e" ,
x"fffdb6",x"fffd5d",x"fffd17",x"fffce5",x"fffcc9",x"fffcc4",x"fffcd6",x"fffcff" ,
x"fffd3c",x"fffd8d",x"fffdef",x"fffe5d",x"fffed6",x"ffff54",x"ffffd4",x"000051" ,
x"0000c9",x"000137",x"000198",x"0001e9",x"000229",x"000256",x"00026f",x"000274" ,
x"000266",x"000247",x"000219",x"0001dd",x"000198",x"00014c",x"0000fe",x"0000af" ,
x"000064",x"000020",x"ffffe5",x"ffffb5",x"ffff92",x"ffff7c",x"ffff74",x"ffff79" ,
x"ffff8a",x"ffffa5",x"ffffc7",x"ffffee",x"000016",x"00003c",x"00005e",x"000077" ,
x"000085",x"000086",x"000078",x"00005a",x"00002c",x"ffffed",x"ffffa1",x"ffff48" ,
x"fffee6",x"fffe7f",x"fffe16",x"fffdb0",x"fffd52",x"fffd01",x"fffcc1",x"fffc97" ,
x"fffc86",x"fffc91",x"fffcbb",x"fffd03",x"fffd6a",x"fffdf0",x"fffe90",x"ffff49" ,
x"000014",x"0000ed",x"0001cd",x"0002ad",x"000385",x"000450",x"000504",x"00059c" ,
x"000611",x"00065f",x"000680",x"000672",x"000635",x"0005c8",x"00052c",x"000466" ,
x"00037b",x"00026f",x"00014c",x"000018",x"fffedd",x"fffda5",x"fffc78",x"fffb61" ,
x"fffa67",x"fff993",x"fff8eb",x"fff875",x"fff835",x"fff82b",x"fff85a",x"fff8bf" ,
x"fff957",x"fffa1d",x"fffb0b",x"fffc19",x"fffd3f",x"fffe73",x"ffffab",x"0000dd" ,
x"000201",x"00030d",x"0003fa",x"0004c0",x"00055c",x"0005c9",x"000605",x"000611" ,
x"0005ef",x"0005a1",x"00052e",x"00049b",x"0003f0",x"000335",x"000272",x"0001af" ,
x"0000f6",x"00004e",x"ffffbc",x"ffff47",x"fffef1",x"fffebe",x"fffead",x"fffebe" ,
x"fffeec",x"ffff33",x"ffff8d",x"fffff3",x"00005d",x"0000c1",x"000117",x"000158" ,
x"00017b",x"00017a",x"000151",x"0000fc",x"00007a",x"ffffcc",x"fffef6",x"fffdfe" ,
x"fffceb",x"fffbc7",x"fffa9e",x"fff97b",x"fff86c",x"fff780",x"fff6c2",x"fff640" ,
x"fff606",x"fff61b",x"fff688",x"fff751",x"fff876",x"fff9f6",x"fffbca",x"fffdea" ,
x"000049",x"0002d7",x"000583",x"000837",x"000adf",x"000d62",x"000faa",x"0011a1" ,
x"001332",x"001449",x"0014d7",x"0014d0",x"00142c",x"0012e6",x"001102",x"000e84" ,
x"000b7a",x"0007f4",x"000407",x"ffffcd",x"fffb62",x"fff6e7",x"fff27c",x"ffee44" ,
x"ffea60",x"ffe6f1",x"ffe416",x"ffe1e8",x"ffe07e",x"ffdfea",x"ffe037",x"ffe169" ,
x"ffe37f",x"ffe670",x"ffea2d",x"ffeea0",x"fff3ae",x"fff935",x"ffff11",x"000518" ,
x"000b20",x"0010fe",x"001685",x"001b8c",x"001fed",x"002384",x"002635",x"0027e8" ,
x"00288d",x"00281c",x"002693",x"0023fb",x"002063",x"001be1",x"001694",x"00109f" ,
x"000a2b",x"000365",x"fffc7d",x"fff5a4",x"ffef0b",x"ffe8e1",x"ffe352",x"ffde86" ,
x"ffda9f",x"ffd7b9",x"ffd5ea",x"07d53e",x"ffd5bb",x"ffd75e",x"ffda1b",x"ffdddd" ,
x"ffe289",x"ffe7fb",x"ffee0d",x"fff491",x"fffb58",x"000230",x"0008ea",x"000f54" ,
x"001542",x"001a8b",x"001f09",x"0022a0",x"002539",x"0026c4",x"00273a",x"00269b" ,
x"0024f0",x"002249",x"001ebd",x"001a6a",x"001572",x"000ffc",x"000a31",x"00043d" ,
x"fffe4b",x"fff886",x"fff317",x"ffee22",x"ffe9c8",x"ffe625",x"ffe34d",x"ffe151" ,
x"ffe039",x"ffe005",x"ffe0b1",x"ffe231",x"ffe474",x"ffe763",x"ffeae3",x"ffeed6" ,
x"fff31c",x"fff792",x"fffc16",x"000087",x"0004c5",x"0008b4",x"000c3a",x"000f41" ,
x"0011ba",x"001399",x"0014d7",x"001572",x"001570",x"0014d7",x"0013b4",x"001218" ,
x"001015",x"000dc0",x"000b31",x"00087e",x"0005bf",x"000308",x"000070",x"fffe08" ,
x"fffbe0",x"fffa04",x"fff87e",x"fff753",x"fff685",x"fff614",x"fff5fa",x"fff632" ,
x"fff6b1",x"fff76c",x"fff858",x"fff965",x"fffa87",x"fffbb0",x"fffcd4",x"fffde7" ,
x"fffee0",x"ffffb6",x"000064",x"0000e6",x"00013c",x"000166",x"000168",x"000145" ,
x"000106",x"0000b0",x"00004d",x"ffffe5",x"ffff80",x"ffff26",x"fffee0",x"fffeb3" ,
x"fffea3",x"fffeb4",x"fffee8",x"ffff3e",x"ffffb3",x"000045",x"0000ed",x"0001a6" ,
x"000268",x"00032b",x"0003e5",x"000490",x"000522",x"000594",x"0005e1",x"000602" ,
x"0005f6",x"0005b9",x"00054b",x"0004b0",x"0003e9",x"0002fd",x"0001f1",x"0000ce" ,
x"ffff9d",x"fffe66",x"fffd34",x"fffc10",x"fffb04",x"fffa19",x"fff955",x"fff8bf" ,
x"fff85d",x"fff831",x"fff83d",x"fff880",x"fff8f9",x"fff9a3",x"fffa78",x"fffb74" ,
x"fffc8c",x"fffdba",x"fffef3",x"00002d",x"000161",x"000284",x"00038e",x"000479" ,
x"00053d",x"0005d7",x"000642",x"00067d",x"000688",x"000665",x"000615",x"00059d" ,
x"000503",x"00044d",x"000381",x"0002a6",x"0001c4",x"0000e3",x"00000a",x"ffff3d" ,
x"fffe85",x"fffde4",x"fffd5e",x"fffcf7",x"fffcaf",x"fffc86",x"fffc7c",x"fffc8e" ,
x"fffcb9",x"fffcfa",x"fffd4c",x"fffdab",x"fffe12",x"fffe7c",x"fffee4",x"ffff47" ,
x"ffffa1",x"ffffee",x"00002d",x"00005d",x"00007b",x"00008a",x"00008a",x"00007c" ,
x"000063",x"000042",x"00001c",x"fffff3",x"ffffcd",x"ffffab",x"ffff90",x"ffff7f" ,
x"ffff7a",x"ffff81",x"ffff97",x"ffffb9",x"ffffe9",x"000023",x"000067",x"0000b1" ,
x"0000ff",x"00014d",x"000198",x"0001dc",x"000217",x"000244",x"000263",x"000270" ,
x"00026a",x"000250",x"000223",x"0001e3",x"000191",x"000130",x"0000c2",x"00004a" ,
x"ffffcd",x"ffff4d",x"fffed0",x"fffe58",x"fffdea",x"fffd8a",x"fffd3a",x"fffcfd" ,
x"fffcd5",x"fffcc4",x"fffcca",x"fffce7",x"fffd1a",x"fffd62",x"fffdbb",x"fffe24" ,
x"fffe99",x"ffff17",x"ffff99",x"00001b",x"00009b",x"000113",x"000181",x"0001e2" ,
x"000232",x"000271",x"00029c",x"0002b4",x"0002b7",x"0002a7",x"000284",x"000251" ,
x"000210",x"0001c3",x"00016e",x"000113",x"0000b5",x"000057",x"fffffd",x"ffffa9" ,
x"ffff5d",x"ffff1b",x"fffee5",x"fffebb",x"fffe9e",x"fffe8f",x"fffe8b",x"fffe94" ,
x"fffea7",x"fffec3",x"fffee5",x"ffff0d",x"ffff38",x"ffff64",x"ffff8f",x"ffffb7" ,
x"ffffdc",x"fffffb",x"000014",x"000027",x"000033",x"000038",x"000037",x"000031" ,
x"000026",x"000018",x"000008",x"fffff8",x"ffffe8",x"ffffda",x"ffffd0",x"ffffc9" ,
x"ffffc8",x"ffffcc",x"ffffd5",x"ffffe4",x"fffff8",x"000010",x"00002c",x"00004a" ,
x"00006a",x"00008a",x"0000a8",x"0000c3",x"0000da",x"0000ec",x"0000f7",x"0000fb" ,
x"0000f8",x"0000ed",x"0000da",x"0000bf",x"00009d",x"000076",x"00004a",x"00001a" ,
x"ffffe8",x"ffffb5",x"ffff83",x"ffff55",x"ffff2a",x"ffff05",x"fffee6",x"fffecf" ,
x"fffec1",x"fffebb",x"fffebf",x"fffecc",x"fffee1",x"fffefd",x"ffff21",x"ffff4b" ,
x"ffff78",x"ffffa9",x"ffffdc",x"00000e",x"00003f",x"00006c",x"000096",x"0000ba" ,
x"0000d8",x"0000ef",x"0000fe",x"000106",x"000106",x"0000ff",x"0000f1",x"0000dd" ,
x"0000c4",x"0000a6",x"000086",x"000063",x"000040",x"00001d",x"fffffc",x"ffffdd" ,
x"ffffc2",x"ffffaa",x"ffff97",x"ffff88",x"ffff7e",x"ffff79",x"ffff79",x"ffff7c" ,
x"ffff84",x"ffff8e",x"ffff9b",x"ffffaa",x"ffffb9",x"ffffc9",x"ffffd9",x"ffffe7" ,
x"fffff4",x"ffffff",x"000007",x"00000e",x"000012",x"000013",x"000012",x"000010" ,
x"00000c",x"000007",x"000001",x"fffffc",x"fffff6",x"fffff2",x"ffffee",x"ffffec" ,
x"ffffec",x"ffffee",x"fffff1",x"fffff6",x"fffffd",x"000006",x"000010",x"00001a" ,
x"000025",x"00002f",x"000039",x"000042",x"00004a",x"000050",x"000053",x"000054" ,
x"000053",x"00004f",x"000048",x"00003f",x"000033",x"000026",x"000017",x"000007" ,
x"fffff6",x"ffffe6",x"ffffd5",x"ffffc6",x"ffffb8",x"ffffad",x"ffffa3",x"ffff9c" ,
x"ffff97",x"ffff96",x"ffff98",x"ffff9c",x"ffffa3",x"ffffad",x"ffffb9",x"ffffc6" ,
x"ffffd5",x"ffffe5",x"fffff5",x"000005",x"000015",x"000024",x"000031",x"00003c" ,
x"000046",x"00004d",x"000052",x"000054",x"000054",x"000051",x"00004d",x"000046" ,
x"00003e",x"000034",x"00002a",x"00001f",x"000013",x"000008",x"fffffe",x"fffff4" ,
x"ffffeb",x"ffffe3",x"ffffdd",x"ffffd8",x"ffffd5",x"ffffd4",x"ffffd3",x"ffffd5" ,
x"ffffd7",x"ffffda",x"ffffdf",x"ffffe3",x"ffffe9",x"ffffee",x"fffff3",x"fffff8" ,
x"fffffc",x"ffffff",x"000002",x"000004",x"000006",x"000006",x"000006",x"000005" ,
x"000004",x"000002",x"000000",x"fffffe",x"fffffc",x"fffffa",x"fffff9",x"fffff8" ,
x"fffff8",x"fffff9",x"fffffa",x"fffffc",x"ffffff",x"000002",x"000006",x"00000a" ,
x"00000f",x"000013",x"000017",x"00001b",x"00001e",x"000021",x"000023",
others=>x"000000"
);
	
	constant COEFFICIENTS_LEN: tCoeffLen := (
		COEFFICIENTS_1_LEN, COEFFICIENTS_2_LEN, COEFFICIENTS_3_LEN, COEFFICIENTS_4_LEN 
		--COEFFICIENTS_5_LEN, COEFFICIENTS_6_LEN, COEFFICIENTS_7_LEN, COEFFICIENTS_8_LEN
	);
	constant COEFFICIENTS: tCoeffArr := (
		COEFFICIENTS_1, COEFFICIENTS_2, COEFFICIENTS_3, COEFFICIENTS_4
		--COEFFICIENTS_5, COEFFICIENTS_6, COEFFICIENTS_7, COEFFICIENTS_8
	);
	
	
	
	
	
	
	
	
	
--	

--	constant COEFFICIENTS: tCoeff := (
--		x"080000",
--		others=>x"000000"
--	);

	

end package constants;